module bitwise_not(out, data);
    input [31:0] data;
    output [31:0] out;

    not NOT0(out[0], data[0]);
    not NOT1(out[1], data[1]);
    not NOT2(out[2], data[2]);
    not NOT3(out[3], data[3]);
    not NOT4(out[4], data[4]);
    not NOT5(out[5], data[5]);
    not NOT6(out[6], data[6]);
    not NOT7(out[7], data[7]);
    not NOT8(out[8], data[8]);
    not NOT9(out[9], data[9]);
    not NOT10(out[10], data[10]);
    not NOT11(out[11], data[11]);
    not NOT12(out[12], data[12]);
    not NOT13(out[13], data[13]);
    not NOT14(out[14], data[14]);
    not NOT15(out[15], data[15]);
    not NOT16(out[16], data[16]);
    not NOT17(out[17], data[17]);
    not NOT18(out[18], data[18]);
    not NOT19(out[19], data[19]);
    not NOT20(out[20], data[20]);
    not NOT21(out[21], data[21]);
    not NOT22(out[22], data[22]);
    not NOT23(out[23], data[23]);
    not NOT24(out[24], data[24]);
    not NOT25(out[25], data[25]);
    not NOT26(out[26], data[26]);
    not NOT27(out[27], data[27]);
    not NOT28(out[28], data[28]);
    not NOT29(out[29], data[29]);
    not NOT30(out[30], data[30]);
    not NOT31(out[31], data[31]);

endmodule